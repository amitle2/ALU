
module NOR2_1 (a,b,c);
 input a;
 input b;
 output c;

 nor nor1 (c,a,b);
endmodule
