
module NOT2_1 (a,b,c);
 input a;
 input b;
 output c;

 not not1 (c,a,b);
endmodule
