
module OR2_1 (a,b,c);
 input a;
 input b;
 output c;

 or or1 (c,a,b);
endmodule
