
module AND2_1 (a,b,c);
 input a;
 input b;
 output c;

 and and1 (c,a,b);
endmodule