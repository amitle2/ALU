
module XOR2_1 (a,b,c);
 input a;
 input b;
 output c;

 xor xor1 (c,a,b);
endmodule
